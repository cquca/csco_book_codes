module disp;
initial begin
$display("\\\t%%\n\"\123");
end
endmodule