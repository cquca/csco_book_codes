always @(a,b)
begin
	e=c&d;
	f=c|d;
end